`include "defines.v"



module ex(
	
	//from id_ex
	input wire[31:0] inst_i,
	input wire[31:0] inst_addr_i,
	input wire[31:0] op1_i,
	input wire[31:0] op2_i,
	input wire[4:0]  rd_addr_i,
	input wire 		 rd_wen_i,
	input wire[31:0] base_addr_i,
	input wire[31:0] offset_addr_i,
	
	//to regs
	output reg[4:0]	 rd_addr_o,
	output reg[31:0] rd_data_o,
	output reg		 rd_wen_o,

	//to ctrl
	output reg[31:0] 	jump_addr_o	,
	output reg 			jump_en_o	,
	output reg 			hold_flag_o	
);

//I type

//extract instructions
	wire[6:0] 	opcode;
	wire[4:0] 	rd;
	wire[2:0] 	func3;
	wire[4:0] 	rs1;
	wire[11:0] 	imm;
	wire[4:0]	rs2;
	wire[6:0]	func7;
	wire[4:0]	shamt;

//I type
	assign opcode 	= inst_i[6:0];
	assign rd 		= inst_i[11:7];
	assign func3 	= inst_i[14:12];
	assign rs1 		= inst_i[19:15];
	assign imm 		= inst_i[31:20];
	assign shamt	= inst_i[24:20];

//R type (others included on top)
	assign rs2 		= inst_i[24:20];
	assign func7	= inst_i[31:25];

// B type
	//wire[31:0]  jump_imm = {{19{inst_i[31]}},inst_i[31], inst_i[7], inst_i[30:25], inst_i[11:8], 1'b0}; //anything infront of bit 13 is all coopied from bit 13, last bit must be 0
	wire		op1_i_equal_op2_i;
	wire		op1_i_less_op2_i_signed;
	wire		op1_i_less_op2_i_unsigned;	

	assign 		op1_i_equal_op2_i			= (op1_i == op2_i)?1'b1:1'b0;
	assign		op1_i_less_op2_i_unsigned 	= (op1_i < op2_i)?1'b1:1'b0;
	assign		op1_i_less_op2_i_signed 	= ($signed (op1_i) < $signed(op2_i))?1'b1:1'b0;

//ALU
	wire[31:0] op1_i_add_op2_i;
	wire[31:0] op1_i_and_op2_i;
	wire[31:0] op1_i_xor_op2_i;
	wire[31:0] op1_i_or_op2_i;
	wire[31:0] op1_i_shift_left_op2_i;
	wire[31:0] op1_i_shift_right_op2_i;
	wire[31:0] base_addr_add_offset_addr;

	assign op1_i_add_op2_i 				= op1_i + op2_i;				//add
	assign op1_i_and_op2_i				= op1_i & op2_i;				//and
	assign op1_i_xor_op2_i				= op1_i ^ op2_i;				//xor
	assign op1_i_or_op2_i				= op1_i | op2_i;				//or
	assign op1_i_shift_left_op2_i		= op1_i << op2_i;				//shift left
	assign op1_i_shift_right_op2_i		= op1_i >> op2_i;				//shift right
	assign base_addr_add_offset_addr	= base_addr_i + offset_addr_i;	//calculate new offset addr

// I Type calculations
	wire[31:0]	SRA_mask;
	assign		SRA_mask = (32'hffff_ffff) >> op2_i [4:0];


	always @(*)begin
		
		case(opcode)

//==================================== I Type ========================================================

			`INST_TYPE_I:begin

				jump_addr_o = 32'b0;
				jump_en_o	= 1'b0;
				hold_flag_o	= 1'b0;

				case(func3)
					
					// ADD IMMEDIATE
					`INST_ADDI:begin
						rd_data_o = op1_i_add_op2_i;
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;
					end

					// SET ON LESS THAN IMMEDIATE
					`INST_SLTI:begin
						rd_data_o = {31'b0, op1_i_less_op2_i_signed};		//tutorial write 30'b0
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;
					end

					// SET ON LESS THAN IMMEDIATE UNISGNED
					`INST_SLTIU:begin
						rd_data_o = {31'b0, op1_i_less_op2_i_unsigned};		//tutorial write 30'b0
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;
					end

					// XOR IMMEDIATE
					`INST_XORI:begin
						rd_data_o = op1_i_xor_op2_i;
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;
					end			

					// OR IMMEDIATE
					`INST_ORI:begin
						rd_data_o = op1_i_or_op2_i;
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;
					end												

					// AND IMMEDIATE
					`INST_ANDI:begin
						rd_data_o = op1_i_and_op2_i;
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;
					end			

					// SHIFT LEFT LOGICAL IMMEDIATE
					`INST_SLLI:begin
						rd_data_o = op1_i_shift_left_op2_i;
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;
					end			

					`INST_SRI: begin
						if(func7[5]== 1'b1) begin 					//SRAI
							rd_data_o = ((op1_i_shift_right_op2_i) & SRA_mask) | (({32{op1_i[31]}}) & ~(SRA_mask));
							rd_addr_o = rd_addr_i;
							rd_wen_o  = 1'b1;							
						end

						else begin									//SRLI
							rd_data_o = op1_i_shift_right_op2_i;
							rd_addr_o = rd_addr_i;
							rd_wen_o  = 1'b1;			
						end
					end					

					default:begin
						rd_data_o = 32'b0;
						rd_addr_o = 5'b0;
						rd_wen_o  = 1'b0;
					end
				endcase
			end

//==================================== R Type ========================================================

			`INST_TYPE_R_M:begin

				jump_addr_o = 32'b0;
				jump_en_o	= 1'b0;
				hold_flag_o	= 1'b0;
									
				case(func3)

					// ADD or SUB
					`INST_ADD_SUB:begin
						if(func7[5] == 1'b0)begin				//ADD
							rd_data_o = op1_i_add_op2_i;
							rd_addr_o = rd_addr_i;
							rd_wen_o  = 1'b1;
						end

						else begin								//SUB
							rd_data_o = op1_i - op2_i;			//rs1-rs2
							rd_addr_o = rd_addr_i;
							rd_wen_o  = 1'b1;
						end
					end

					// SHIFT LEFT LOGICAL
					`INST_SLL:begin

						rd_data_o = op1_i_shift_left_op2_i;		//After 4 bit no point
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;

					end

					// SET LESS THAN
					`INST_SLT:begin

						rd_data_o = {31'b0, op1_i_less_op2_i_signed};		
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;

					end

					// SET LESS THAN UNSIGNED
					`INST_SLTU:begin

						rd_data_o = {31'b0, op1_i_less_op2_i_unsigned};	
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;

					end

					// XOR
					`INST_XOR:begin

						rd_data_o = op1_i_xor_op2_i;		
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;

					end

					// OR
					`INST_OR:begin

						rd_data_o = op1_i_or_op2_i;		
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;

					end

					// AND
					`INST_AND:begin

						rd_data_o = op1_i_and_op2_i;		
						rd_addr_o = rd_addr_i;
						rd_wen_o  = 1'b1;

					end

					// SHIFT RIGHT
					`INST_SR:begin

						if(func7[5]== 1'b1) begin 					//SRA
							rd_data_o = ((op1_i_shift_right_op2_i) & SRA_mask) | (({32{op1_i[31]}}) & ~(SRA_mask));
							rd_addr_o = rd_addr_i;
							rd_wen_o  = 1'b1;							
						end

						else begin									//SRL
							rd_data_o = op1_i_shift_right_op2_i;
							rd_addr_o = rd_addr_i;
							rd_wen_o  = 1'b1;			
						end

					end

					default:begin
						rd_data_o = 32'b0;
						rd_addr_o = 5'b0;
						rd_wen_o  = 1'b0;
					end
				endcase
			end	

//==================================== B Type ========================================================

			`INST_TYPE_B:begin
				rd_data_o = 32'b0;
				rd_addr_o = 5'b0;
				rd_wen_o  = 1'b0;
				case(func3)

					// BRANCH EQUAL
					`INST_BEQ:begin
						jump_addr_o = base_addr_add_offset_addr;
						jump_en_o	= op1_i_equal_op2_i;		//EQUAL, JUMP
						hold_flag_o	= 1'b0;			
					end					

					// BRANCH NOT EQUAL
					`INST_BNE:begin
						jump_addr_o = base_addr_add_offset_addr;
						jump_en_o	= ~op1_i_equal_op2_i;		//NOT EQUAL, JUMP
						hold_flag_o	= 1'b0;					
					end

					// BRANCH LESS THAN
					`INST_BLT:begin
						jump_addr_o = base_addr_add_offset_addr;
						jump_en_o	= op1_i_less_op2_i_signed;		//LESS THAN, JUMP
						hold_flag_o	= 1'b0;					
					end

					//BRANCH GREATER THAN
					`INST_BGE:begin
						jump_addr_o = base_addr_add_offset_addr;
						jump_en_o	= ~op1_i_less_op2_i_signed;		//GREATER THAN, JUMP
						hold_flag_o	= 1'b0;					
					end

					// BRANCH LESS THAN UNSIGNED
					`INST_BLTU:begin
						jump_addr_o = base_addr_add_offset_addr;
						jump_en_o	= op1_i_less_op2_i_unsigned;			//LESS THAN(UNSIGNED), JUMP
						hold_flag_o	= 1'b0;					
					end

					// BRANCH GREATER THAN UNSIGNED
					`INST_BGEU:begin
						jump_addr_o = base_addr_add_offset_addr;
						jump_en_o	= ~op1_i_less_op2_i_unsigned;			//GREATER THAN (UNSIGNED), JUMP
						hold_flag_o	= 1'b0;					
					end

					default:begin
						jump_addr_o = 32'b0;
						jump_en_o	= 1'b0;
						hold_flag_o	= 1'b0;	
					end
				endcase
			end

//==================================== J Type ========================================================

			`INST_JAL:begin
				rd_data_o = op1_i_add_op2_i;
				rd_addr_o = rd_addr_i;
				rd_wen_o  = 1'b1;
				jump_addr_o = base_addr_add_offset_addr;
				jump_en_o	= 1'b1;
				hold_flag_o	= 1'b0;	
			end

			`INST_JALR:begin
				rd_data_o = op1_i_add_op2_i;
				rd_addr_o = rd_addr_i;
				rd_wen_o  = 1'b1;
				jump_addr_o = base_addr_add_offset_addr;
				jump_en_o	= 1'b1;
				hold_flag_o	= 1'b0;	
			end

//==================================== U Type ========================================================

			`INST_LUI:begin
				rd_data_o 	= op1_i;
				rd_addr_o 	= rd_addr_i;
				rd_wen_o  	= 1'b1;
				jump_addr_o = 32'b0;
				jump_en_o	= 1'b0;
				hold_flag_o	= 1'b0;	
			end					

			`INST_AUIPC:begin
				rd_data_o 	= op1_i_add_op2_i;
				rd_addr_o 	= rd_addr_i;
				rd_wen_o  	= 1'b1;
				jump_addr_o = 32'b0;
				jump_en_o	= 1'b0;
				hold_flag_o	= 1'b0;	
			end		

			default:begin
				rd_data_o = 32'b0;
				rd_addr_o = 5'b0;
				rd_wen_o  = 1'b0;
				jump_addr_o = 32'b0;
				jump_en_o	= 1'b0;
				hold_flag_o	= 1'b0;	
			end
		endcase
	
	end

endmodule